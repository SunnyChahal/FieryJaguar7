module card7seg (SW, HEX0);

input [3:0] SW;
output [6:0] HEX0;
		
   // Your code for Phase 2 goes here.  Be sure to check the Slide Set 2 notes,
   // since one of the slides almost gives away the answer here.  I wrote this as
   // a single combinational always block containing a single case statement, but 
   // there are other ways to do it.
	
endmodule
