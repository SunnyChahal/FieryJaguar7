module reg4 (in, load, rst, clk, out) begin
	input [3:0] in;
	input load, rst, clk;
	output [3:0] out;
	
	//always block for a 4-bit wide register with asynchronous reset
	
endmodule